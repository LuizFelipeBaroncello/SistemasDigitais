library verilog;
use verilog.vl_types.all;
entity topoPart4_vlg_vec_tst is
end topoPart4_vlg_vec_tst;
