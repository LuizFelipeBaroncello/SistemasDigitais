library verilog;
use verilog.vl_types.all;
entity part2 is
    port(
        Clk             : in     vl_logic;
        D               : in     vl_logic;
        Q               : out    vl_logic;
        QN              : out    vl_logic
    );
end part2;
